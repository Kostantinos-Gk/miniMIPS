--MIPS Part_6
--MemoryInstruction_MIPS
--Memory Set specialy for the implementation of FINAL_PROJECT
--27/05/2020, Konstantinos Gkousaris, 711171073, UniWA

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;


ENTITY instrMemoryMIPS IS PORT (
		Addr : IN STD_LOGIC_VECTOR(3 downto 0);
		C : out STD_LOGIC_VECTOR(31 downto 0));
END instrMemoryMIPS;

ARCHITECTURE behavioral OF instrMemoryMIPS IS

TYPE rom16x32 IS ARRAY (0 TO 15) OF STD_LOGIC_VECTOR(31 downto 0);
       
        --give default 
	SIGNAL instrmem : rom16x32 := (    			--Instruction Set
		"00000000010001100010000000100000",		--add $4 $2 $6
		"00000000010001100010100000100010",		--sub $5 $2 $6
		"00000000000000000000000000000000",		
		"00000000000000000000000000000000",		
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 		 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",             
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111");
BEGIN
	C <= instrmem(to_integer(unsigned(Addr)));

END;