--MIPS Part_4
--MemoryInstruction
--27/05/2020, Konstantinos Gkousaris, 711171073, UniWA

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;


ENTITY instrMemory IS PORT (
		Addr : IN STD_LOGIC_VECTOR(3 downto 0);
		C : out STD_LOGIC_VECTOR(31 downto 0));
END instrMemory;

ARCHITECTURE arch1 OF instrMemory IS

TYPE rom16x32 IS ARRAY (0 TO 15) OF STD_LOGIC_VECTOR(31 downto 0);
       
        --give default 
	SIGNAL instrmem : rom16x32 := (    			--Instruction Set
		"00000001001010000101000000100010",		--sub  $5, $1, $0
		"00000001001010000101000000100100",		--and  $5, $4, $3
		"00000000101001100010000000100000",		--add $4, $5, $6 
		"00000000100000010000000000000000",		--jump to address 0
		"11111111111111111111111111111111",
		"00000000000000000000000000000000", 		 
		"11111111111111111111111111111111",
		"00000000100000010000000000000000",             
		"11111111111111111111111111111111",
		"00000000101001100010000000100000",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111");
BEGIN
	C <= instrmem(to_integer(unsigned(Addr)));

END arch1;